module top.v(

);
endmodule