module test_bench(

);